---------------------------------------------------------------------------------- 
-- Create Date: 06/04/2025 04:16:55 PM
-- Design Name: 
-- Module Name: Control_Unit - Behavioral
-- Project Name: 
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity Control_Unit is
  Port (
       -- IR 
       D : in std_logic;
       ld: in std_logic
       
   );
end Control_Unit;

architecture Behavioral of Control_Unit is

begin


end Behavioral;
